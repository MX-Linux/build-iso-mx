   1)  Standard
   2)  automount       Montera enheter automatiskt när de pluggas in
   3)  noautomount     Stäng av all extra montering och automontering
