   1)  Standard
   2)  checkmd5        Kontrollera live-mediums integritet
   3)  checkfs         Kontrollera LiveUSB och persistens ext2/3/4 filsystem
   4)  toram           Kopiera det komprimerade filsystemet till RAM
   5)  i915_invert     Invert video on some Intel graphics systems
   6)  no_i915_invert  Disable Intel graphics invert
   7)  from=usb        Slutför start från en LiveUSB
   8)  from=hd         Slutför start från en hårddisk
   9)  hwclock=ask     Få hjälp av systemet att avgöra klockans inställning
  10)  hwclock=utc     Hårdvaru-klockan använder UTC (Endast Linuxsystem)
  11)  hwclock=local   Hårdvaru-klocka använder lokal tid (Windows system)
  12)  password        Ändra lösenord före start
  13)  nostore         Stäng av LiveUSB-lagringsfunktionen (Endast LiveUSB)
  14)  dostore         Använd LiveUSB-lagringsfunktionen (Endast LiveUSB)
  15)  savestate       Spara en del filer vid omstarter (Endast LiveUSB)
  16)  nosavestate     Spara inte filer vid omstarter (Endast LiveUSB)
