   1)  Standard
   2)  persist_all     Spara root i RAM, spara home på disken (spara root vid avstängning)
   3)  persist_root    Spara root och home i RAM sedan sparade vid avstängning
   4)  persist_static  Spara root och home på disken med home separat på disken
   5)  p_static_root   Spara root och home på disken tillsammans
   6)  persist_home    Bara home-persistens
   7)  frugal_persist  Frugal med root i RAM och home på disken
   8)  frugal_root     Frugal med root och home i RAM sedan sparade vid avstängning
   9)  frugal_static   Frugal med root på disken och home separat på disken
  10)  f_static_root   Frugal med root och home på disken tillsammans
  11)  frugal_home     Frugal med endast home-persistens
  12)  frugal_only     Bara Frugal, ingen persistens
